module and1(input D0, input D1,output wire SelData);
       assign SelData = D0 & D1;
endmodule