module instructionmemory(addr, instruction);
    
   //input reset;
	input [31:0] addr;
	output reg [31:0] instruction;
	reg [31:0] Imem [31:0];
	
	integer i;
	wire [29:0] shifted_addr;
	assign shifted_addr= addr[31:2];

	initial begin
        //Imem[1] <= 32'b0000000_01010_00000_000_00100_0010011;   //      ADDI x4, x0, 10 
		  
      Imem[0] <= 32'h0000_0000;
      //Imem[1] <= 32'h00200193;   // addi x2, x0, 1
      Imem[2] <= 32'h00100193;  // addi x3, x0, 1
      Imem[3] <= 32'h00600293;//  addi x5, x0, 6
      Imem[4] <= 32'h00020233; // add x4, x4, x0
      Imem[5] <= 32'h00218133; //  add x2, x3, x2
      Imem[6] <= 32'h000103b3;  // add x7, x2, x0
      Imem[7] <= 32'h00018133; //add x2, x3, x0
      Imem[8] <= 32'h000381b3;   // add x3, x7, x0 
      Imem[9] <= 32'h00120213; //  addi x4, x4, 1
      Imem[10] <= 32'hfe428de3;// beq x5, x4, -6

		  Imem[1] <= 32'h01088933;   //      add x18 , x17, x16
		  //Imem[2] <= 32'h0108e9b3;    //     or x19 , x17, x16
		  //Imem[2] <= 32'h01060633;  // add x12, x12, x16
		  //Imem[3] <= 32'h01060633;  // add x12, x12, x16
        //Imem[2] <= 32'h00962223;   //      sw x9, 4(x0)
		  //Imem[3] <= 32'h0108ca33;   //      xor x20 , x17, x16
        //Imem[4] <= 32'h00542503;		//     lw x10, 5(x8)
        //Imem[2] <= 32'h0108e9b3;   //     or x19 , x17, x16
        //Imem[3] <= 32'h0108ca33;   //      xor x20 , x17, x16 
		  //Imem[4]  <= 32'h01181463; // bne x16, x17, 8
		  //Imem[5] <= 32'h01180263; // beq x16, x17, 4
       // Imem[6] <= 32'h3e860713;   //      addi x14, x12, 1000
        //Imem[7] <= 32'h3e85c513;   //      xori x10, x11, 1000                                                                                     
        //Imem[6] <= 32'b1111111_00000_00101_000_10001_1100011;   //      BEQ x5, x0, Sort 
        //Imem[7] <= 32'b0000000_00000_00101_010_00111_0000011;   //      LW x7, 0(x5)        
        //Imem[8] <= 32'b0000000_00000_00110_010_01000_0000011;   //      LW x8, 0(x6)        
        //Imem[9] <= 32'b0000000_00111_01000_010_01001_0110011;   //      SLT x9, x8, x7      
        //Imem[10] <= 32'b0000000_00000_01001_001_01100_1100011;   //      BNE x9, x0                                                                                      
        Imem[11] <= 32'b0000000_01000_00101_010_00000_0100011;   //      SW x8, 0(x5)        
        Imem[12] <= 32'b0000000_00111_00110_010_00000_0100011;   //      SW x7, 0(x6)                            
        Imem[13] <= 32'b1111111_11100_00101_000_00101_0010011;   //      ADDI x5, x5, -4     
        Imem[14] <= 32'b1111111_11100_00101_000_00110_0010011;   //      ADDI x6, x5, -4     
        Imem[15] <= 32'b1111110_11101_11111_111_01010_1101111;   //      JAL x10, Itr      
        Imem[16] <= 32'b0000000_00000_00000_010_00001_0000011;   //      LW x1, 0(x0)
        Imem[17] <= 32'b0000000_00100_00000_010_00010_0000011;   //      LW x2, 4(x0)
        Imem[18] <= 32'b0000000_01000_00000_010_00011_0000011;   //      LW x3, 8(x0)
        Imem[19] <= 32'b0000000_01100_00000_010_00100_0000011;   //      LW x4, 12(x0)
        Imem[20] <= 32'b0000000_10000_00000_010_00101_0000011;   //      LW x5, 16(x0)
        Imem[21] <= 32'b0000000_10100_00000_010_00110_0000011;   //      LW x6, 20(x0)
        Imem[22] <= 32'b0000000_11000_00000_010_00111_0000011;   //      LW x7, 24(x0)
        Imem[23] <= 32'b0000000_11100_00000_010_01000_0000011;   //      LW x8, 28(x0)
        Imem[24] <= 32'b0000001_00000_00000_010_01001_0000011;   //      LW x9, 32(x0)
        Imem[25] <= 32'b0000001_00100_00000_010_01010_0000011;   //      LW x10, 36(x0)
        
	     for (i = 26; i < 31; i = i + 1) begin
            Imem[i] = 32'h0000_0000;
        end
    end
    
  always@(*)begin
    instruction = Imem[shifted_addr];
  end


endmodule