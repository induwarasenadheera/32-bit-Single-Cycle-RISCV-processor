module processor();


endmodule
